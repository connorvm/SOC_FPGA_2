-- Authors: Connor Van Meter & Alex Salois
-- EELE 468
-- HW_4

library IEEE;
use IEEE.numeric_std.all;
use IEEE.std_logic_1164.all;

entity yo_block is

  generic (W_bits   : positive;
           F_bits   : positive);

  port (clock   : in std_logic;
  	    reset   : in std_logic;
	      y_in    : in  unsigned(W_bits - 1 downto 0);
 	      x	      : in  unsigned(W_bits - 1 downto 0);
	      out_n   : out unsigned(W_bits - 1 downto 0));
end entity;

architecture yo_block_arch of yo_block is

  signal y_relay_0 : unsigned(W_bits - 1 downto 0) := (others => '0');
  signal y_relay_1 : unsigned(W_bits - 1 downto 0) := (others => '0');
  signal y_relay_2 : unsigned(W_bits - 1 downto 0) := (others => '0');
  signal y_relay_3 : unsigned(W_bits - 1 downto 0) := (others => '0');
  signal x_relay_0 : unsigned(W_bits - 1 downto 0) := (others => '0');
  signal Y_next    : unsigned(4*W_bits - 1 downto 0) := (others => '0');
  signal xy_square : unsigned(3*W_bits - 1 downto 0) := (others => '0');
  signal minus     : unsigned(3*W_bits - 1 downto 0) := (others => '0');
  signal square    : unsigned(2*W_bits - 1 downto 0) := (others => '0');
  signal top	     : unsigned(4*W_bits - 1 downto 0) := (others => '0');

  constant three : unsigned(3*W_bits - 1 downto 0) := (3*F_bits + 1 downto 3*F_bits => '1', others => '0');

  begin
    --y_(n+1) = (y_n(3 -x(y_n)^2))/2
  process (clock, reset)
  begin
    if(reset = '0') then
	out_n <= "0";
    elsif(rising_edge(clock)) then
    	square 	  <= y_in * y_in; -- square y_current
    	xy_square <= x_relay_0 * square;
	    minus 	  <= three - xy_square;
	    top       <= y_relay_3 * minus;
      y_next 	  <= shift_right(top, 1); -- divide by 2
    	out_n 	<= y_next((4*F_bits -1) + (W_bits - F_bits) downto 4*F_bits -  F_bits);

    end if;
  end process;

  process (clock, reset)
  begin
    if(reset = '0') then
	--out_n <= "0";
    elsif(rising_edge(clock)) then
      y_relay_0 <= y_in;
	    y_relay_1 <= y_relay_0;
	    y_relay_2 <= y_relay_1;
	    y_relay_3 <= y_relay_2;
	    x_relay_0 <= x;

    end if;
  end process;

end architecture;